module converter_onecold_bin (

)
endmodule